magic
tech sky130A
magscale 1 2
timestamp 1647626135
<< nwell >>
rect -40 -62 235 563
<< nsubdiff >>
rect 68 275 162 299
rect 68 241 98 275
rect 135 241 162 275
rect 68 207 162 241
rect 68 173 98 207
rect 135 173 162 207
rect 68 144 162 173
<< nsubdiffcont >>
rect 98 241 135 275
rect 98 173 135 207
<< poly >>
rect -40 405 235 435
rect -9 22 21 405
rect 63 32 147 48
rect 63 22 79 32
rect -40 -8 79 22
rect 63 -20 79 -8
rect 131 22 147 32
rect 190 22 220 405
rect 131 -8 235 22
rect 131 -20 147 -8
rect 63 -36 147 -20
<< polycont >>
rect 79 -20 131 32
<< locali >>
rect 39 275 190 299
rect 39 273 98 275
rect 39 239 42 273
rect 76 241 98 273
rect 135 241 190 275
rect 76 239 190 241
rect 39 207 190 239
rect 39 190 98 207
rect 39 156 42 190
rect 76 173 98 190
rect 135 173 190 207
rect 76 156 190 173
rect 39 152 190 156
rect 63 32 147 48
rect 63 -20 79 32
rect 131 -20 147 32
rect 63 -36 147 -20
<< viali >>
rect 42 239 76 273
rect 42 156 76 190
rect 79 -20 131 32
<< metal1 >>
rect 13 299 41 563
rect 13 273 82 299
rect 172 276 200 563
rect 13 239 42 273
rect 76 239 82 273
rect 13 190 82 239
rect 13 156 42 190
rect 76 156 82 190
rect 13 144 82 156
rect 144 152 200 276
rect 13 -62 41 144
rect 69 32 144 46
rect 69 -20 79 32
rect 131 -20 144 32
rect 69 -34 144 -20
rect 172 -62 200 152
<< via1 >>
rect 79 -20 131 32
<< metal2 >>
rect -40 276 235 316
rect -40 193 235 226
rect -40 80 235 118
rect 73 32 137 80
rect 73 -20 79 32
rect 131 -20 137 32
rect 73 -27 137 -20
<< properties >>
string FIXED_BBOX @z���
<< end >>
