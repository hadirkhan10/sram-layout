magic
tech sky130A
magscale 1 2
timestamp 1647626531
<< pwell >>
rect -24 -32 251 593
<< psubdiff >>
rect 84 307 178 329
rect 84 273 112 307
rect 149 273 178 307
rect 84 239 178 273
rect 84 205 111 239
rect 148 205 178 239
rect 84 174 178 205
<< psubdiffcont >>
rect 112 273 149 307
rect 111 205 148 239
<< poly >>
rect -24 435 251 465
rect 7 52 38 435
rect 80 62 164 79
rect 80 52 96 62
rect -24 22 96 52
rect 80 10 96 22
rect 148 52 164 62
rect 206 52 236 435
rect 148 22 251 52
rect 148 10 164 22
rect 80 -5 164 10
<< polycont >>
rect 96 10 148 62
<< locali >>
rect 56 308 207 329
rect 56 307 176 308
rect 56 273 112 307
rect 149 274 176 307
rect 149 273 207 274
rect 56 239 207 273
rect 56 205 111 239
rect 148 236 207 239
rect 148 205 174 236
rect 56 202 174 205
rect 56 182 207 202
rect 80 62 164 79
rect 80 10 96 62
rect 148 10 164 62
rect 80 -5 164 10
<< viali >>
rect 176 274 210 308
rect 174 202 208 236
rect 96 10 148 62
<< metal1 >>
rect 29 329 57 593
rect 188 329 216 593
rect 29 174 84 329
rect 147 308 216 329
rect 147 274 176 308
rect 210 274 216 308
rect 147 236 216 274
rect 147 202 174 236
rect 208 202 216 236
rect 147 174 216 202
rect 29 -32 57 174
rect 85 62 160 77
rect 85 10 96 62
rect 148 10 160 62
rect 85 -3 160 10
rect 188 -32 216 174
<< via1 >>
rect 96 10 148 62
<< metal2 >>
rect -24 306 251 346
rect -24 223 251 256
rect -24 110 251 148
rect 90 62 154 110
rect 90 10 96 62
rect 148 10 154 62
rect 90 4 154 10
<< end >>
