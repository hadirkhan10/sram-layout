magic
tech sky130A
magscale 1 2
timestamp 1647626135
<< nwell >>
rect 148 -365 408 260
<< pwell >>
rect -124 -365 65 260
<< scnmos >>
rect -12 102 60 132
rect -12 -63 60 -33
rect -12 -159 60 -129
rect -12 -311 60 -281
<< pmos >>
rect 184 -63 268 -27
rect 184 -165 268 -129
<< ndiff >>
rect -12 195 60 205
rect -12 161 6 195
rect 40 161 60 195
rect -12 132 60 161
rect -12 59 60 102
rect -12 25 9 59
rect 43 25 60 59
rect -12 -33 60 25
rect -118 -78 -66 -70
rect -12 -78 60 -63
rect -124 -79 60 -78
rect -124 -113 -108 -79
rect -74 -113 60 -79
rect -124 -114 60 -113
rect -118 -122 -66 -114
rect -12 -129 60 -114
rect -12 -224 60 -159
rect -12 -258 5 -224
rect 39 -258 60 -224
rect -12 -281 60 -258
rect -12 -323 60 -311
rect -12 -357 6 -323
rect 40 -357 60 -323
rect -12 -365 60 -357
<< pdiff >>
rect 184 60 268 83
rect 184 26 211 60
rect 245 26 268 60
rect 184 -27 268 26
rect 184 -83 268 -63
rect 322 -79 372 -67
rect 322 -83 330 -79
rect 184 -113 330 -83
rect 364 -113 372 -79
rect 184 -129 268 -113
rect 322 -125 372 -113
rect 184 -224 268 -165
rect 184 -258 209 -224
rect 243 -258 268 -224
rect 184 -266 268 -258
<< ndiffc >>
rect 6 161 40 195
rect 9 25 43 59
rect -108 -113 -74 -79
rect 5 -258 39 -224
rect 6 -357 40 -323
<< pdiffc >>
rect 211 26 245 60
rect 330 -113 364 -79
rect 209 -258 243 -224
<< poly >>
rect -124 102 -12 132
rect 60 102 408 132
rect 84 -27 153 -17
rect 84 -28 184 -27
rect 84 -33 103 -28
rect -38 -63 -12 -33
rect 60 -62 103 -33
rect 137 -62 184 -28
rect 60 -63 184 -62
rect 268 -63 294 -27
rect 84 -72 150 -63
rect 82 -124 151 -114
rect 82 -129 98 -124
rect -38 -159 -12 -129
rect 60 -158 98 -129
rect 132 -129 151 -124
rect 132 -158 184 -129
rect 60 -159 184 -158
rect 82 -165 184 -159
rect 268 -165 296 -129
rect 82 -169 151 -165
rect -124 -311 -12 -281
rect 60 -311 408 -281
<< polycont >>
rect 103 -62 137 -28
rect 98 -158 132 -124
<< locali >>
rect -12 192 6 195
rect -22 161 6 192
rect 40 192 60 195
rect 40 161 80 192
rect -22 158 80 161
rect 136 158 285 192
rect -7 59 211 60
rect -7 25 9 59
rect 43 26 211 59
rect 245 26 268 60
rect 43 25 268 26
rect -7 22 268 25
rect 84 -28 150 -12
rect 84 -29 103 -28
rect 5 -62 103 -29
rect 137 -62 150 -28
rect 5 -63 150 -62
rect -124 -79 -54 -78
rect -124 -113 -108 -79
rect -74 -113 -54 -79
rect -124 -114 -54 -113
rect 5 -221 45 -63
rect 84 -78 150 -63
rect 82 -124 148 -112
rect 82 -158 98 -124
rect 132 -125 148 -124
rect 202 -125 236 22
rect 132 -158 236 -125
rect 319 -79 380 -63
rect 319 -113 330 -79
rect 364 -113 380 -79
rect 319 -129 380 -113
rect 82 -159 236 -158
rect 82 -176 148 -159
rect -11 -224 269 -221
rect -11 -258 5 -224
rect 39 -258 209 -224
rect 243 -258 269 -224
rect -21 -357 6 -323
rect 40 -357 171 -323
rect 227 -357 286 -323
rect 6 -361 40 -357
<< viali >>
rect 80 158 136 192
rect -108 -113 -74 -79
rect 330 -113 364 -79
rect 171 -357 227 -323
<< metal1 >>
rect -124 -55 -69 260
rect 86 199 131 260
rect 68 192 150 199
rect 68 158 80 192
rect 136 158 150 192
rect 68 146 150 158
rect -124 -61 -50 -55
rect -124 -113 -108 -61
rect -56 -113 -50 -61
rect -124 -119 -50 -113
rect -124 -122 -67 -119
rect -124 -365 -69 -122
rect 86 -365 131 146
rect 180 -315 215 260
rect 332 31 408 260
rect 322 25 408 31
rect 322 -27 328 25
rect 380 -27 408 25
rect 322 -33 408 -27
rect 328 -63 408 -33
rect 323 -79 408 -63
rect 323 -113 330 -79
rect 364 -113 408 -79
rect 323 -125 408 -113
rect 159 -323 241 -315
rect 159 -357 171 -323
rect 227 -357 241 -323
rect 159 -365 241 -357
rect 332 -365 408 -125
<< via1 >>
rect -108 -79 -56 -61
rect -108 -113 -74 -79
rect -74 -113 -56 -79
rect 328 -27 380 25
<< metal2 >>
rect 322 25 386 31
rect 322 13 328 25
rect -124 -27 328 13
rect 380 13 386 25
rect 380 -27 408 13
rect 322 -33 386 -27
rect -114 -61 -50 -55
rect -114 -77 -108 -61
rect -124 -110 -108 -77
rect -114 -113 -108 -110
rect -56 -77 -50 -61
rect -56 -110 408 -77
rect -56 -113 -50 -110
rect -114 -119 -50 -113
rect -124 -223 408 -185
<< labels >>
rlabel pwell -65 -357 -53 -343 1 VNB
port 1 n
rlabel metal1 -93 -348 -74 -329 1 VGND
port 2 n
rlabel metal1 96 66 115 85 1 BL
port 3 n
rlabel metal1 187 66 206 85 1 BR
port 4 n
rlabel poly 141 107 160 126 1 WL
port 5 n
rlabel poly 135 -308 154 -289 1 WL
port 5 n
rlabel nwell 377 -350 400 -326 1 VPB
port 6 n
rlabel metal1 337 -349 360 -325 1 VPWR
port 7 n
<< end >>
